library IEEE;
 use IEEE.std_logic_1164.all;
 
 entity RxUnit is
   port (
     clk, reset       : in  std_logic;
     enable           : in  std_logic;
     read             : in  std_logic;
     rxd              : in  std_logic;
     data             : out std_logic_vector(7 downto 0);
     Ferr, OErr, DRdy : out std_logic);
 end RxUnit;
 
 architecture RxUnit_arch of RxUnit is
 begin
     data <= "00000000";
     Ferr <= '0';
     OErr <= '0';
     DRdy <= '0';
 end RxUnit_arch;
